MACRO FIVE_TRANSISTOR_OTA
  ORIGIN 0 0 ;
  FOREIGN FIVE_TRANSISTOR_OTA 0 0 ;
  SIZE 28.51 BY 35.03 ;
  PIN ID
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 14.05 2.78 14.33 7.3 ;
    END
  END ID
  PIN VOUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 13.19 14.12 13.47 20.32 ;
      LAYER M3 ;
        RECT 13.62 21.68 13.9 27.88 ;
      LAYER M3 ;
        RECT 13.19 19.975 13.47 20.345 ;
      LAYER M4 ;
        RECT 13.33 19.76 13.76 20.56 ;
      LAYER M3 ;
        RECT 13.62 20.16 13.9 21.84 ;
    END
  END VOUT
  PIN VINP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 13.62 10.34 13.9 16.54 ;
    END
  END VINP
  PIN VINN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 14.05 9.92 14.33 16.12 ;
    END
  END VINN
  OBS 
  LAYER M2 ;
        RECT 1.98 6.58 22.96 6.86 ;
  LAYER M3 ;
        RECT 14.48 13.7 14.76 19.9 ;
  LAYER M2 ;
        RECT 14.46 6.58 14.78 6.86 ;
  LAYER M3 ;
        RECT 14.48 6.72 14.76 13.86 ;
  LAYER M2 ;
        RECT 14.46 6.58 14.78 6.86 ;
  LAYER M3 ;
        RECT 14.48 6.56 14.76 6.88 ;
  LAYER M2 ;
        RECT 14.46 6.58 14.78 6.86 ;
  LAYER M3 ;
        RECT 14.48 6.56 14.76 6.88 ;
  LAYER M3 ;
        RECT 12.76 14.54 13.04 20.74 ;
  LAYER M3 ;
        RECT 13.19 21.26 13.47 31.66 ;
  LAYER M3 ;
        RECT 12.76 20.58 13.04 21 ;
  LAYER M2 ;
        RECT 12.9 20.86 13.33 21.14 ;
  LAYER M3 ;
        RECT 13.19 21 13.47 21.42 ;
  LAYER M2 ;
        RECT 12.74 20.86 13.06 21.14 ;
  LAYER M3 ;
        RECT 12.76 20.84 13.04 21.16 ;
  LAYER M2 ;
        RECT 13.17 20.86 13.49 21.14 ;
  LAYER M3 ;
        RECT 13.19 20.84 13.47 21.16 ;
  LAYER M2 ;
        RECT 12.74 20.86 13.06 21.14 ;
  LAYER M3 ;
        RECT 12.76 20.84 13.04 21.16 ;
  LAYER M2 ;
        RECT 13.17 20.86 13.49 21.14 ;
  LAYER M3 ;
        RECT 13.19 20.84 13.47 21.16 ;
  LAYER M1 ;
        RECT 25.245 3.695 25.495 7.225 ;
  LAYER M1 ;
        RECT 25.245 2.435 25.495 3.445 ;
  LAYER M1 ;
        RECT 25.245 0.335 25.495 1.345 ;
  LAYER M1 ;
        RECT 26.535 3.695 26.785 7.225 ;
  LAYER M1 ;
        RECT 23.955 3.695 24.205 7.225 ;
  LAYER M1 ;
        RECT 22.665 3.695 22.915 7.225 ;
  LAYER M1 ;
        RECT 22.665 2.435 22.915 3.445 ;
  LAYER M1 ;
        RECT 22.665 0.335 22.915 1.345 ;
  LAYER M1 ;
        RECT 21.375 3.695 21.625 7.225 ;
  LAYER M1 ;
        RECT 20.085 3.695 20.335 7.225 ;
  LAYER M1 ;
        RECT 20.085 2.435 20.335 3.445 ;
  LAYER M1 ;
        RECT 20.085 0.335 20.335 1.345 ;
  LAYER M1 ;
        RECT 18.795 3.695 19.045 7.225 ;
  LAYER M1 ;
        RECT 17.505 3.695 17.755 7.225 ;
  LAYER M1 ;
        RECT 17.505 2.435 17.755 3.445 ;
  LAYER M1 ;
        RECT 17.505 0.335 17.755 1.345 ;
  LAYER M1 ;
        RECT 16.215 3.695 16.465 7.225 ;
  LAYER M1 ;
        RECT 14.925 3.695 15.175 7.225 ;
  LAYER M1 ;
        RECT 14.925 2.435 15.175 3.445 ;
  LAYER M1 ;
        RECT 14.925 0.335 15.175 1.345 ;
  LAYER M1 ;
        RECT 13.635 3.695 13.885 7.225 ;
  LAYER M1 ;
        RECT 12.345 3.695 12.595 7.225 ;
  LAYER M1 ;
        RECT 12.345 2.435 12.595 3.445 ;
  LAYER M1 ;
        RECT 12.345 0.335 12.595 1.345 ;
  LAYER M1 ;
        RECT 11.055 3.695 11.305 7.225 ;
  LAYER M1 ;
        RECT 9.765 3.695 10.015 7.225 ;
  LAYER M1 ;
        RECT 9.765 2.435 10.015 3.445 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 1.345 ;
  LAYER M1 ;
        RECT 8.475 3.695 8.725 7.225 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.185 2.435 7.435 3.445 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 1.345 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M1 ;
        RECT 4.605 3.695 4.855 7.225 ;
  LAYER M1 ;
        RECT 4.605 2.435 4.855 3.445 ;
  LAYER M1 ;
        RECT 4.605 0.335 4.855 1.345 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M1 ;
        RECT 2.025 3.695 2.275 7.225 ;
  LAYER M1 ;
        RECT 2.025 2.435 2.275 3.445 ;
  LAYER M1 ;
        RECT 2.025 0.335 2.275 1.345 ;
  LAYER M1 ;
        RECT 0.735 3.695 0.985 7.225 ;
  LAYER M2 ;
        RECT 1.98 2.8 25.54 3.08 ;
  LAYER M2 ;
        RECT 4.56 7 25.54 7.28 ;
  LAYER M2 ;
        RECT 0.69 6.16 26.83 6.44 ;
  LAYER M2 ;
        RECT 1.98 0.7 25.54 0.98 ;
  LAYER M3 ;
        RECT 14.05 2.78 14.33 7.3 ;
  LAYER M2 ;
        RECT 1.98 6.58 22.96 6.86 ;
  LAYER M3 ;
        RECT 13.19 0.68 13.47 6.46 ;
  LAYER M1 ;
        RECT 2.025 21.335 2.275 24.865 ;
  LAYER M1 ;
        RECT 2.025 25.115 2.275 26.125 ;
  LAYER M1 ;
        RECT 2.025 27.215 2.275 30.745 ;
  LAYER M1 ;
        RECT 2.025 30.995 2.275 32.005 ;
  LAYER M1 ;
        RECT 2.025 33.095 2.275 34.105 ;
  LAYER M1 ;
        RECT 0.735 21.335 0.985 24.865 ;
  LAYER M1 ;
        RECT 0.735 27.215 0.985 30.745 ;
  LAYER M1 ;
        RECT 3.315 21.335 3.565 24.865 ;
  LAYER M1 ;
        RECT 3.315 27.215 3.565 30.745 ;
  LAYER M1 ;
        RECT 4.605 21.335 4.855 24.865 ;
  LAYER M1 ;
        RECT 4.605 25.115 4.855 26.125 ;
  LAYER M1 ;
        RECT 4.605 27.215 4.855 30.745 ;
  LAYER M1 ;
        RECT 4.605 30.995 4.855 32.005 ;
  LAYER M1 ;
        RECT 4.605 33.095 4.855 34.105 ;
  LAYER M1 ;
        RECT 5.895 21.335 6.145 24.865 ;
  LAYER M1 ;
        RECT 5.895 27.215 6.145 30.745 ;
  LAYER M1 ;
        RECT 7.185 21.335 7.435 24.865 ;
  LAYER M1 ;
        RECT 7.185 25.115 7.435 26.125 ;
  LAYER M1 ;
        RECT 7.185 27.215 7.435 30.745 ;
  LAYER M1 ;
        RECT 7.185 30.995 7.435 32.005 ;
  LAYER M1 ;
        RECT 7.185 33.095 7.435 34.105 ;
  LAYER M1 ;
        RECT 8.475 21.335 8.725 24.865 ;
  LAYER M1 ;
        RECT 8.475 27.215 8.725 30.745 ;
  LAYER M1 ;
        RECT 9.765 21.335 10.015 24.865 ;
  LAYER M1 ;
        RECT 9.765 25.115 10.015 26.125 ;
  LAYER M1 ;
        RECT 9.765 27.215 10.015 30.745 ;
  LAYER M1 ;
        RECT 9.765 30.995 10.015 32.005 ;
  LAYER M1 ;
        RECT 9.765 33.095 10.015 34.105 ;
  LAYER M1 ;
        RECT 11.055 21.335 11.305 24.865 ;
  LAYER M1 ;
        RECT 11.055 27.215 11.305 30.745 ;
  LAYER M1 ;
        RECT 12.345 21.335 12.595 24.865 ;
  LAYER M1 ;
        RECT 12.345 25.115 12.595 26.125 ;
  LAYER M1 ;
        RECT 12.345 27.215 12.595 30.745 ;
  LAYER M1 ;
        RECT 12.345 30.995 12.595 32.005 ;
  LAYER M1 ;
        RECT 12.345 33.095 12.595 34.105 ;
  LAYER M1 ;
        RECT 13.635 21.335 13.885 24.865 ;
  LAYER M1 ;
        RECT 13.635 27.215 13.885 30.745 ;
  LAYER M1 ;
        RECT 14.925 21.335 15.175 24.865 ;
  LAYER M1 ;
        RECT 14.925 25.115 15.175 26.125 ;
  LAYER M1 ;
        RECT 14.925 27.215 15.175 30.745 ;
  LAYER M1 ;
        RECT 14.925 30.995 15.175 32.005 ;
  LAYER M1 ;
        RECT 14.925 33.095 15.175 34.105 ;
  LAYER M1 ;
        RECT 16.215 21.335 16.465 24.865 ;
  LAYER M1 ;
        RECT 16.215 27.215 16.465 30.745 ;
  LAYER M1 ;
        RECT 17.505 21.335 17.755 24.865 ;
  LAYER M1 ;
        RECT 17.505 25.115 17.755 26.125 ;
  LAYER M1 ;
        RECT 17.505 27.215 17.755 30.745 ;
  LAYER M1 ;
        RECT 17.505 30.995 17.755 32.005 ;
  LAYER M1 ;
        RECT 17.505 33.095 17.755 34.105 ;
  LAYER M1 ;
        RECT 18.795 21.335 19.045 24.865 ;
  LAYER M1 ;
        RECT 18.795 27.215 19.045 30.745 ;
  LAYER M1 ;
        RECT 20.085 21.335 20.335 24.865 ;
  LAYER M1 ;
        RECT 20.085 25.115 20.335 26.125 ;
  LAYER M1 ;
        RECT 20.085 27.215 20.335 30.745 ;
  LAYER M1 ;
        RECT 20.085 30.995 20.335 32.005 ;
  LAYER M1 ;
        RECT 20.085 33.095 20.335 34.105 ;
  LAYER M1 ;
        RECT 21.375 21.335 21.625 24.865 ;
  LAYER M1 ;
        RECT 21.375 27.215 21.625 30.745 ;
  LAYER M1 ;
        RECT 22.665 21.335 22.915 24.865 ;
  LAYER M1 ;
        RECT 22.665 25.115 22.915 26.125 ;
  LAYER M1 ;
        RECT 22.665 27.215 22.915 30.745 ;
  LAYER M1 ;
        RECT 22.665 30.995 22.915 32.005 ;
  LAYER M1 ;
        RECT 22.665 33.095 22.915 34.105 ;
  LAYER M1 ;
        RECT 23.955 21.335 24.205 24.865 ;
  LAYER M1 ;
        RECT 23.955 27.215 24.205 30.745 ;
  LAYER M1 ;
        RECT 25.245 21.335 25.495 24.865 ;
  LAYER M1 ;
        RECT 25.245 25.115 25.495 26.125 ;
  LAYER M1 ;
        RECT 25.245 27.215 25.495 30.745 ;
  LAYER M1 ;
        RECT 25.245 30.995 25.495 32.005 ;
  LAYER M1 ;
        RECT 25.245 33.095 25.495 34.105 ;
  LAYER M1 ;
        RECT 26.535 21.335 26.785 24.865 ;
  LAYER M1 ;
        RECT 26.535 27.215 26.785 30.745 ;
  LAYER M2 ;
        RECT 1.98 25.48 25.54 25.76 ;
  LAYER M2 ;
        RECT 1.98 21.28 22.96 21.56 ;
  LAYER M2 ;
        RECT 4.56 21.7 25.54 21.98 ;
  LAYER M2 ;
        RECT 0.69 22.12 26.83 22.4 ;
  LAYER M2 ;
        RECT 1.98 31.36 25.54 31.64 ;
  LAYER M2 ;
        RECT 4.56 27.16 25.54 27.44 ;
  LAYER M2 ;
        RECT 1.98 27.58 22.96 27.86 ;
  LAYER M2 ;
        RECT 0.69 28 26.83 28.28 ;
  LAYER M2 ;
        RECT 1.98 33.46 25.54 33.74 ;
  LAYER M3 ;
        RECT 13.19 21.26 13.47 31.66 ;
  LAYER M3 ;
        RECT 13.62 21.68 13.9 27.88 ;
  LAYER M3 ;
        RECT 14.05 22.1 14.33 33.76 ;
  LAYER M1 ;
        RECT 2.025 17.135 2.275 20.665 ;
  LAYER M1 ;
        RECT 2.025 15.875 2.275 16.885 ;
  LAYER M1 ;
        RECT 2.025 11.255 2.275 14.785 ;
  LAYER M1 ;
        RECT 2.025 9.995 2.275 11.005 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 8.905 ;
  LAYER M1 ;
        RECT 0.735 17.135 0.985 20.665 ;
  LAYER M1 ;
        RECT 0.735 11.255 0.985 14.785 ;
  LAYER M1 ;
        RECT 3.315 17.135 3.565 20.665 ;
  LAYER M1 ;
        RECT 3.315 11.255 3.565 14.785 ;
  LAYER M1 ;
        RECT 4.605 17.135 4.855 20.665 ;
  LAYER M1 ;
        RECT 4.605 15.875 4.855 16.885 ;
  LAYER M1 ;
        RECT 4.605 11.255 4.855 14.785 ;
  LAYER M1 ;
        RECT 4.605 9.995 4.855 11.005 ;
  LAYER M1 ;
        RECT 4.605 7.895 4.855 8.905 ;
  LAYER M1 ;
        RECT 5.895 17.135 6.145 20.665 ;
  LAYER M1 ;
        RECT 5.895 11.255 6.145 14.785 ;
  LAYER M1 ;
        RECT 7.185 17.135 7.435 20.665 ;
  LAYER M1 ;
        RECT 7.185 15.875 7.435 16.885 ;
  LAYER M1 ;
        RECT 7.185 11.255 7.435 14.785 ;
  LAYER M1 ;
        RECT 7.185 9.995 7.435 11.005 ;
  LAYER M1 ;
        RECT 7.185 7.895 7.435 8.905 ;
  LAYER M1 ;
        RECT 8.475 17.135 8.725 20.665 ;
  LAYER M1 ;
        RECT 8.475 11.255 8.725 14.785 ;
  LAYER M1 ;
        RECT 9.765 17.135 10.015 20.665 ;
  LAYER M1 ;
        RECT 9.765 15.875 10.015 16.885 ;
  LAYER M1 ;
        RECT 9.765 11.255 10.015 14.785 ;
  LAYER M1 ;
        RECT 9.765 9.995 10.015 11.005 ;
  LAYER M1 ;
        RECT 9.765 7.895 10.015 8.905 ;
  LAYER M1 ;
        RECT 11.055 17.135 11.305 20.665 ;
  LAYER M1 ;
        RECT 11.055 11.255 11.305 14.785 ;
  LAYER M1 ;
        RECT 12.345 17.135 12.595 20.665 ;
  LAYER M1 ;
        RECT 12.345 15.875 12.595 16.885 ;
  LAYER M1 ;
        RECT 12.345 11.255 12.595 14.785 ;
  LAYER M1 ;
        RECT 12.345 9.995 12.595 11.005 ;
  LAYER M1 ;
        RECT 12.345 7.895 12.595 8.905 ;
  LAYER M1 ;
        RECT 13.635 17.135 13.885 20.665 ;
  LAYER M1 ;
        RECT 13.635 11.255 13.885 14.785 ;
  LAYER M1 ;
        RECT 14.925 17.135 15.175 20.665 ;
  LAYER M1 ;
        RECT 14.925 15.875 15.175 16.885 ;
  LAYER M1 ;
        RECT 14.925 11.255 15.175 14.785 ;
  LAYER M1 ;
        RECT 14.925 9.995 15.175 11.005 ;
  LAYER M1 ;
        RECT 14.925 7.895 15.175 8.905 ;
  LAYER M1 ;
        RECT 16.215 17.135 16.465 20.665 ;
  LAYER M1 ;
        RECT 16.215 11.255 16.465 14.785 ;
  LAYER M1 ;
        RECT 17.505 17.135 17.755 20.665 ;
  LAYER M1 ;
        RECT 17.505 15.875 17.755 16.885 ;
  LAYER M1 ;
        RECT 17.505 11.255 17.755 14.785 ;
  LAYER M1 ;
        RECT 17.505 9.995 17.755 11.005 ;
  LAYER M1 ;
        RECT 17.505 7.895 17.755 8.905 ;
  LAYER M1 ;
        RECT 18.795 17.135 19.045 20.665 ;
  LAYER M1 ;
        RECT 18.795 11.255 19.045 14.785 ;
  LAYER M1 ;
        RECT 20.085 17.135 20.335 20.665 ;
  LAYER M1 ;
        RECT 20.085 15.875 20.335 16.885 ;
  LAYER M1 ;
        RECT 20.085 11.255 20.335 14.785 ;
  LAYER M1 ;
        RECT 20.085 9.995 20.335 11.005 ;
  LAYER M1 ;
        RECT 20.085 7.895 20.335 8.905 ;
  LAYER M1 ;
        RECT 21.375 17.135 21.625 20.665 ;
  LAYER M1 ;
        RECT 21.375 11.255 21.625 14.785 ;
  LAYER M1 ;
        RECT 22.665 17.135 22.915 20.665 ;
  LAYER M1 ;
        RECT 22.665 15.875 22.915 16.885 ;
  LAYER M1 ;
        RECT 22.665 11.255 22.915 14.785 ;
  LAYER M1 ;
        RECT 22.665 9.995 22.915 11.005 ;
  LAYER M1 ;
        RECT 22.665 7.895 22.915 8.905 ;
  LAYER M1 ;
        RECT 23.955 17.135 24.205 20.665 ;
  LAYER M1 ;
        RECT 23.955 11.255 24.205 14.785 ;
  LAYER M1 ;
        RECT 25.245 17.135 25.495 20.665 ;
  LAYER M1 ;
        RECT 25.245 15.875 25.495 16.885 ;
  LAYER M1 ;
        RECT 25.245 11.255 25.495 14.785 ;
  LAYER M1 ;
        RECT 25.245 9.995 25.495 11.005 ;
  LAYER M1 ;
        RECT 25.245 7.895 25.495 8.905 ;
  LAYER M1 ;
        RECT 26.535 17.135 26.785 20.665 ;
  LAYER M1 ;
        RECT 26.535 11.255 26.785 14.785 ;
  LAYER M2 ;
        RECT 1.98 20.44 22.96 20.72 ;
  LAYER M2 ;
        RECT 4.56 20.02 25.54 20.3 ;
  LAYER M2 ;
        RECT 1.98 16.24 22.96 16.52 ;
  LAYER M2 ;
        RECT 4.56 15.82 25.54 16.1 ;
  LAYER M2 ;
        RECT 0.69 19.6 26.83 19.88 ;
  LAYER M2 ;
        RECT 4.56 14.56 25.54 14.84 ;
  LAYER M2 ;
        RECT 1.98 14.14 22.96 14.42 ;
  LAYER M2 ;
        RECT 4.56 10.36 25.54 10.64 ;
  LAYER M2 ;
        RECT 1.98 9.94 22.96 10.22 ;
  LAYER M2 ;
        RECT 0.69 13.72 26.83 14 ;
  LAYER M2 ;
        RECT 1.98 8.26 25.54 8.54 ;
  LAYER M3 ;
        RECT 12.76 14.54 13.04 20.74 ;
  LAYER M3 ;
        RECT 13.19 14.12 13.47 20.32 ;
  LAYER M3 ;
        RECT 13.62 10.34 13.9 16.54 ;
  LAYER M3 ;
        RECT 14.05 9.92 14.33 16.12 ;
  LAYER M3 ;
        RECT 14.48 13.7 14.76 19.9 ;
  END 
END FIVE_TRANSISTOR_OTA
