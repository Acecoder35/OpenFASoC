MACRO BUFFER
  ORIGIN 0 0 ;
  FOREIGN BUFFER 0 0 ;
  SIZE 12.04 BY 15.12 ;
  PIN VSS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 3.3 0.68 3.58 6.88 ;
      LAYER M3 ;
        RECT 8.46 0.68 8.74 6.88 ;
      LAYER M3 ;
        RECT 3.3 1.075 3.58 1.445 ;
      LAYER M2 ;
        RECT 3.44 1.12 8.6 1.4 ;
      LAYER M3 ;
        RECT 8.46 1.075 8.74 1.445 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 3.3 8.24 3.58 14.44 ;
      LAYER M3 ;
        RECT 8.46 8.24 8.74 14.44 ;
      LAYER M3 ;
        RECT 3.3 8.635 3.58 9.005 ;
      LAYER M2 ;
        RECT 3.44 8.68 8.6 8.96 ;
      LAYER M3 ;
        RECT 8.46 8.635 8.74 9.005 ;
    END
  END VDD
  PIN IN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 7.14 2.8 10.92 3.08 ;
      LAYER M2 ;
        RECT 7.14 12.04 10.92 12.32 ;
      LAYER M2 ;
        RECT 7.58 2.8 7.9 3.08 ;
      LAYER M3 ;
        RECT 7.6 2.94 7.88 12.18 ;
      LAYER M2 ;
        RECT 7.58 12.04 7.9 12.32 ;
    END
  END IN
  PIN OUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.12 7 4.9 7.28 ;
      LAYER M2 ;
        RECT 1.12 7.84 4.9 8.12 ;
      LAYER M2 ;
        RECT 1.56 7 1.88 7.28 ;
      LAYER M3 ;
        RECT 1.58 7.14 1.86 7.98 ;
      LAYER M2 ;
        RECT 1.56 7.84 1.88 8.12 ;
    END
  END OUT
  OBS 
  LAYER M2 ;
        RECT 1.12 2.8 4.9 3.08 ;
  LAYER M2 ;
        RECT 1.12 12.04 4.9 12.32 ;
  LAYER M2 ;
        RECT 7.14 7 10.92 7.28 ;
  LAYER M2 ;
        RECT 7.14 7.84 10.92 8.12 ;
  LAYER M2 ;
        RECT 1.13 2.8 1.45 3.08 ;
  LAYER M3 ;
        RECT 1.15 2.94 1.43 12.18 ;
  LAYER M2 ;
        RECT 1.13 12.04 1.45 12.32 ;
  LAYER M2 ;
        RECT 4.73 2.8 6.45 3.08 ;
  LAYER M1 ;
        RECT 6.325 2.94 6.575 7.14 ;
  LAYER M2 ;
        RECT 6.45 7 7.31 7.28 ;
  LAYER M2 ;
        RECT 7.15 7 7.47 7.28 ;
  LAYER M3 ;
        RECT 7.17 7.14 7.45 7.98 ;
  LAYER M2 ;
        RECT 7.15 7.84 7.47 8.12 ;
  LAYER M2 ;
        RECT 1.13 2.8 1.45 3.08 ;
  LAYER M3 ;
        RECT 1.15 2.78 1.43 3.1 ;
  LAYER M2 ;
        RECT 1.13 12.04 1.45 12.32 ;
  LAYER M3 ;
        RECT 1.15 12.02 1.43 12.34 ;
  LAYER M2 ;
        RECT 1.13 2.8 1.45 3.08 ;
  LAYER M3 ;
        RECT 1.15 2.78 1.43 3.1 ;
  LAYER M2 ;
        RECT 1.13 12.04 1.45 12.32 ;
  LAYER M3 ;
        RECT 1.15 12.02 1.43 12.34 ;
  LAYER M1 ;
        RECT 6.325 2.855 6.575 3.025 ;
  LAYER M2 ;
        RECT 6.28 2.8 6.62 3.08 ;
  LAYER M1 ;
        RECT 6.325 7.055 6.575 7.225 ;
  LAYER M2 ;
        RECT 6.28 7 6.62 7.28 ;
  LAYER M2 ;
        RECT 1.13 2.8 1.45 3.08 ;
  LAYER M3 ;
        RECT 1.15 2.78 1.43 3.1 ;
  LAYER M2 ;
        RECT 1.13 12.04 1.45 12.32 ;
  LAYER M3 ;
        RECT 1.15 12.02 1.43 12.34 ;
  LAYER M1 ;
        RECT 6.325 2.855 6.575 3.025 ;
  LAYER M2 ;
        RECT 6.28 2.8 6.62 3.08 ;
  LAYER M1 ;
        RECT 6.325 7.055 6.575 7.225 ;
  LAYER M2 ;
        RECT 6.28 7 6.62 7.28 ;
  LAYER M2 ;
        RECT 1.13 2.8 1.45 3.08 ;
  LAYER M3 ;
        RECT 1.15 2.78 1.43 3.1 ;
  LAYER M2 ;
        RECT 1.13 12.04 1.45 12.32 ;
  LAYER M3 ;
        RECT 1.15 12.02 1.43 12.34 ;
  LAYER M1 ;
        RECT 6.325 2.855 6.575 3.025 ;
  LAYER M2 ;
        RECT 6.28 2.8 6.62 3.08 ;
  LAYER M1 ;
        RECT 6.325 7.055 6.575 7.225 ;
  LAYER M2 ;
        RECT 6.28 7 6.62 7.28 ;
  LAYER M2 ;
        RECT 1.13 2.8 1.45 3.08 ;
  LAYER M3 ;
        RECT 1.15 2.78 1.43 3.1 ;
  LAYER M2 ;
        RECT 1.13 12.04 1.45 12.32 ;
  LAYER M3 ;
        RECT 1.15 12.02 1.43 12.34 ;
  LAYER M2 ;
        RECT 7.15 7 7.47 7.28 ;
  LAYER M3 ;
        RECT 7.17 6.98 7.45 7.3 ;
  LAYER M2 ;
        RECT 7.15 7.84 7.47 8.12 ;
  LAYER M3 ;
        RECT 7.17 7.82 7.45 8.14 ;
  LAYER M1 ;
        RECT 6.325 2.855 6.575 3.025 ;
  LAYER M2 ;
        RECT 6.28 2.8 6.62 3.08 ;
  LAYER M1 ;
        RECT 6.325 7.055 6.575 7.225 ;
  LAYER M2 ;
        RECT 6.28 7 6.62 7.28 ;
  LAYER M2 ;
        RECT 1.13 2.8 1.45 3.08 ;
  LAYER M3 ;
        RECT 1.15 2.78 1.43 3.1 ;
  LAYER M2 ;
        RECT 1.13 12.04 1.45 12.32 ;
  LAYER M3 ;
        RECT 1.15 12.02 1.43 12.34 ;
  LAYER M2 ;
        RECT 7.15 7 7.47 7.28 ;
  LAYER M3 ;
        RECT 7.17 6.98 7.45 7.3 ;
  LAYER M2 ;
        RECT 7.15 7.84 7.47 8.12 ;
  LAYER M3 ;
        RECT 7.17 7.82 7.45 8.14 ;
  LAYER M1 ;
        RECT 10.625 3.695 10.875 7.225 ;
  LAYER M1 ;
        RECT 10.625 2.435 10.875 3.445 ;
  LAYER M1 ;
        RECT 10.625 0.335 10.875 1.345 ;
  LAYER M1 ;
        RECT 11.055 3.695 11.305 7.225 ;
  LAYER M1 ;
        RECT 10.195 3.695 10.445 7.225 ;
  LAYER M1 ;
        RECT 9.765 3.695 10.015 7.225 ;
  LAYER M1 ;
        RECT 9.765 2.435 10.015 3.445 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 1.345 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M1 ;
        RECT 8.905 3.695 9.155 7.225 ;
  LAYER M1 ;
        RECT 8.905 2.435 9.155 3.445 ;
  LAYER M1 ;
        RECT 8.905 0.335 9.155 1.345 ;
  LAYER M1 ;
        RECT 8.475 3.695 8.725 7.225 ;
  LAYER M1 ;
        RECT 8.045 3.695 8.295 7.225 ;
  LAYER M1 ;
        RECT 8.045 2.435 8.295 3.445 ;
  LAYER M1 ;
        RECT 8.045 0.335 8.295 1.345 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.185 2.435 7.435 3.445 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 1.345 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M2 ;
        RECT 7.14 0.7 10.92 0.98 ;
  LAYER M2 ;
        RECT 6.71 6.58 11.35 6.86 ;
  LAYER M2 ;
        RECT 7.14 7 10.92 7.28 ;
  LAYER M2 ;
        RECT 7.14 2.8 10.92 3.08 ;
  LAYER M3 ;
        RECT 8.46 0.68 8.74 6.88 ;
  LAYER M1 ;
        RECT 1.165 3.695 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.165 2.435 1.415 3.445 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 1.345 ;
  LAYER M1 ;
        RECT 0.735 3.695 0.985 7.225 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M1 ;
        RECT 2.025 3.695 2.275 7.225 ;
  LAYER M1 ;
        RECT 2.025 2.435 2.275 3.445 ;
  LAYER M1 ;
        RECT 2.025 0.335 2.275 1.345 ;
  LAYER M1 ;
        RECT 2.455 3.695 2.705 7.225 ;
  LAYER M1 ;
        RECT 2.885 3.695 3.135 7.225 ;
  LAYER M1 ;
        RECT 2.885 2.435 3.135 3.445 ;
  LAYER M1 ;
        RECT 2.885 0.335 3.135 1.345 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.745 2.435 3.995 3.445 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 1.345 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M1 ;
        RECT 4.605 3.695 4.855 7.225 ;
  LAYER M1 ;
        RECT 4.605 2.435 4.855 3.445 ;
  LAYER M1 ;
        RECT 4.605 0.335 4.855 1.345 ;
  LAYER M1 ;
        RECT 5.035 3.695 5.285 7.225 ;
  LAYER M2 ;
        RECT 1.12 0.7 4.9 0.98 ;
  LAYER M2 ;
        RECT 0.69 6.58 5.33 6.86 ;
  LAYER M2 ;
        RECT 1.12 7 4.9 7.28 ;
  LAYER M2 ;
        RECT 1.12 2.8 4.9 3.08 ;
  LAYER M3 ;
        RECT 3.3 0.68 3.58 6.88 ;
  LAYER M1 ;
        RECT 10.625 7.895 10.875 11.425 ;
  LAYER M1 ;
        RECT 10.625 11.675 10.875 12.685 ;
  LAYER M1 ;
        RECT 10.625 13.775 10.875 14.785 ;
  LAYER M1 ;
        RECT 11.055 7.895 11.305 11.425 ;
  LAYER M1 ;
        RECT 10.195 7.895 10.445 11.425 ;
  LAYER M1 ;
        RECT 9.765 7.895 10.015 11.425 ;
  LAYER M1 ;
        RECT 9.765 11.675 10.015 12.685 ;
  LAYER M1 ;
        RECT 9.765 13.775 10.015 14.785 ;
  LAYER M1 ;
        RECT 9.335 7.895 9.585 11.425 ;
  LAYER M1 ;
        RECT 8.905 7.895 9.155 11.425 ;
  LAYER M1 ;
        RECT 8.905 11.675 9.155 12.685 ;
  LAYER M1 ;
        RECT 8.905 13.775 9.155 14.785 ;
  LAYER M1 ;
        RECT 8.475 7.895 8.725 11.425 ;
  LAYER M1 ;
        RECT 8.045 7.895 8.295 11.425 ;
  LAYER M1 ;
        RECT 8.045 11.675 8.295 12.685 ;
  LAYER M1 ;
        RECT 8.045 13.775 8.295 14.785 ;
  LAYER M1 ;
        RECT 7.615 7.895 7.865 11.425 ;
  LAYER M1 ;
        RECT 7.185 7.895 7.435 11.425 ;
  LAYER M1 ;
        RECT 7.185 11.675 7.435 12.685 ;
  LAYER M1 ;
        RECT 7.185 13.775 7.435 14.785 ;
  LAYER M1 ;
        RECT 6.755 7.895 7.005 11.425 ;
  LAYER M2 ;
        RECT 7.14 14.14 10.92 14.42 ;
  LAYER M2 ;
        RECT 6.71 8.26 11.35 8.54 ;
  LAYER M2 ;
        RECT 7.14 7.84 10.92 8.12 ;
  LAYER M2 ;
        RECT 7.14 12.04 10.92 12.32 ;
  LAYER M3 ;
        RECT 8.46 8.24 8.74 14.44 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 14.785 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 11.425 ;
  LAYER M1 ;
        RECT 2.025 11.675 2.275 12.685 ;
  LAYER M1 ;
        RECT 2.025 13.775 2.275 14.785 ;
  LAYER M1 ;
        RECT 2.455 7.895 2.705 11.425 ;
  LAYER M1 ;
        RECT 2.885 7.895 3.135 11.425 ;
  LAYER M1 ;
        RECT 2.885 11.675 3.135 12.685 ;
  LAYER M1 ;
        RECT 2.885 13.775 3.135 14.785 ;
  LAYER M1 ;
        RECT 3.315 7.895 3.565 11.425 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 11.425 ;
  LAYER M1 ;
        RECT 3.745 11.675 3.995 12.685 ;
  LAYER M1 ;
        RECT 3.745 13.775 3.995 14.785 ;
  LAYER M1 ;
        RECT 4.175 7.895 4.425 11.425 ;
  LAYER M1 ;
        RECT 4.605 7.895 4.855 11.425 ;
  LAYER M1 ;
        RECT 4.605 11.675 4.855 12.685 ;
  LAYER M1 ;
        RECT 4.605 13.775 4.855 14.785 ;
  LAYER M1 ;
        RECT 5.035 7.895 5.285 11.425 ;
  LAYER M2 ;
        RECT 1.12 14.14 4.9 14.42 ;
  LAYER M2 ;
        RECT 0.69 8.26 5.33 8.54 ;
  LAYER M2 ;
        RECT 1.12 7.84 4.9 8.12 ;
  LAYER M2 ;
        RECT 1.12 12.04 4.9 12.32 ;
  LAYER M3 ;
        RECT 3.3 8.24 3.58 14.44 ;
  END 
END BUFFER
