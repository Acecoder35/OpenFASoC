MACRO CP
  ORIGIN 0 0 ;
  FOREIGN CP 0 0 ;
  SIZE 11.18 BY 22.68 ;
  PIN VSS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 1.58 8.24 1.86 14.44 ;
      LAYER M3 ;
        RECT 9.32 8.24 9.6 14.44 ;
      LAYER M3 ;
        RECT 8.03 15.8 8.31 22 ;
      LAYER M3 ;
        RECT 5.02 16.22 5.3 22 ;
      LAYER M3 ;
        RECT 1.58 8.635 1.86 9.005 ;
      LAYER M2 ;
        RECT 1.72 8.68 9.46 8.96 ;
      LAYER M3 ;
        RECT 9.32 8.635 9.6 9.005 ;
      LAYER M3 ;
        RECT 9.32 14.28 9.6 15.12 ;
      LAYER M2 ;
        RECT 8.17 14.98 9.46 15.26 ;
      LAYER M3 ;
        RECT 8.03 15.12 8.31 15.96 ;
      LAYER M3 ;
        RECT 8.03 16.615 8.31 16.985 ;
      LAYER M2 ;
        RECT 5.16 16.66 8.17 16.94 ;
      LAYER M3 ;
        RECT 5.02 16.615 5.3 16.985 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 1.58 0.68 1.86 6.88 ;
      LAYER M3 ;
        RECT 4.59 1.1 4.87 6.88 ;
      LAYER M3 ;
        RECT 9.32 0.68 9.6 6.88 ;
      LAYER M3 ;
        RECT 2.87 15.8 3.15 22 ;
      LAYER M3 ;
        RECT 1.58 1.495 1.86 1.865 ;
      LAYER M2 ;
        RECT 1.72 1.54 4.73 1.82 ;
      LAYER M3 ;
        RECT 4.59 1.495 4.87 1.865 ;
      LAYER M3 ;
        RECT 4.59 1.915 4.87 2.285 ;
      LAYER M2 ;
        RECT 4.73 1.96 9.46 2.24 ;
      LAYER M3 ;
        RECT 9.32 1.915 9.6 2.285 ;
      LAYER M3 ;
        RECT 1.58 6.72 1.86 7.56 ;
      LAYER M2 ;
        RECT 1.72 7.42 3.01 7.7 ;
      LAYER M3 ;
        RECT 2.87 7.56 3.15 15.96 ;
    END
  END VDD
  PIN UP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.26 7 1.46 7.28 ;
      LAYER M2 ;
        RECT 0.26 7.84 1.46 8.12 ;
      LAYER M2 ;
        RECT 0.27 7 0.59 7.28 ;
      LAYER M1 ;
        RECT 0.305 7.14 0.555 7.98 ;
      LAYER M2 ;
        RECT 0.27 7.84 0.59 8.12 ;
      LAYER M2 ;
        RECT 3.7 9.94 4.9 10.22 ;
      LAYER M2 ;
        RECT 1.29 7.84 3.44 8.12 ;
      LAYER M1 ;
        RECT 3.315 7.98 3.565 10.08 ;
      LAYER M2 ;
        RECT 3.44 9.94 3.87 10.22 ;
    END
  END UP
  PIN DN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 9.72 7 10.92 7.28 ;
      LAYER M2 ;
        RECT 9.72 7.84 10.92 8.12 ;
      LAYER M2 ;
        RECT 10.59 7 10.91 7.28 ;
      LAYER M1 ;
        RECT 10.625 7.14 10.875 7.98 ;
      LAYER M2 ;
        RECT 10.59 7.84 10.91 8.12 ;
      LAYER M2 ;
        RECT 7.14 10.36 8.34 10.64 ;
      LAYER M2 ;
        RECT 8.17 7.84 9.89 8.12 ;
      LAYER M1 ;
        RECT 8.045 7.98 8.295 10.5 ;
      LAYER M2 ;
        RECT 8.01 10.36 8.33 10.64 ;
    END
  END DN
  PIN OUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 7.14 7 8.34 7.28 ;
      LAYER M2 ;
        RECT 3.7 14.14 4.9 14.42 ;
      LAYER M2 ;
        RECT 5.59 7 7.31 7.28 ;
      LAYER M1 ;
        RECT 5.465 7.14 5.715 14.28 ;
      LAYER M2 ;
        RECT 4.73 14.14 5.59 14.42 ;
    END
  END OUT
  OBS 
  LAYER M3 ;
        RECT 5.88 15.38 6.16 19.9 ;
  LAYER M3 ;
        RECT 5.02 8.24 5.3 14.02 ;
  LAYER M2 ;
        RECT 4.99 15.82 6.19 16.1 ;
  LAYER M3 ;
        RECT 5.02 13.86 5.3 15.12 ;
  LAYER M2 ;
        RECT 5.16 14.98 5.59 15.26 ;
  LAYER M3 ;
        RECT 5.45 15.12 5.73 15.96 ;
  LAYER M2 ;
        RECT 5.43 15.82 5.75 16.1 ;
  LAYER M2 ;
        RECT 5 14.98 5.32 15.26 ;
  LAYER M3 ;
        RECT 5.02 14.96 5.3 15.28 ;
  LAYER M2 ;
        RECT 5.43 14.98 5.75 15.26 ;
  LAYER M3 ;
        RECT 5.45 14.96 5.73 15.28 ;
  LAYER M2 ;
        RECT 5.43 15.82 5.75 16.1 ;
  LAYER M3 ;
        RECT 5.45 15.8 5.73 16.12 ;
  LAYER M2 ;
        RECT 5 14.98 5.32 15.26 ;
  LAYER M3 ;
        RECT 5.02 14.96 5.3 15.28 ;
  LAYER M2 ;
        RECT 5.43 14.98 5.75 15.26 ;
  LAYER M3 ;
        RECT 5.45 14.96 5.73 15.28 ;
  LAYER M2 ;
        RECT 5.43 15.82 5.75 16.1 ;
  LAYER M3 ;
        RECT 5.45 15.8 5.73 16.12 ;
  LAYER M3 ;
        RECT 3.73 0.26 4.01 4.78 ;
  LAYER M2 ;
        RECT 3.7 0.7 4.9 0.98 ;
  LAYER M3 ;
        RECT 6.74 0.68 7.02 6.88 ;
  LAYER M3 ;
        RECT 6.74 8.24 7.02 14.44 ;
  LAYER M2 ;
        RECT 4.73 0.7 6.02 0.98 ;
  LAYER M3 ;
        RECT 5.88 0.84 6.16 1.26 ;
  LAYER M2 ;
        RECT 6.02 1.12 6.88 1.4 ;
  LAYER M3 ;
        RECT 6.74 1.075 7.02 1.445 ;
  LAYER M3 ;
        RECT 6.74 6.72 7.02 8.4 ;
  LAYER M2 ;
        RECT 5.86 0.7 6.18 0.98 ;
  LAYER M3 ;
        RECT 5.88 0.68 6.16 1 ;
  LAYER M2 ;
        RECT 5.86 1.12 6.18 1.4 ;
  LAYER M3 ;
        RECT 5.88 1.1 6.16 1.42 ;
  LAYER M2 ;
        RECT 6.72 1.12 7.04 1.4 ;
  LAYER M3 ;
        RECT 6.74 1.1 7.02 1.42 ;
  LAYER M2 ;
        RECT 5.86 0.7 6.18 0.98 ;
  LAYER M3 ;
        RECT 5.88 0.68 6.16 1 ;
  LAYER M2 ;
        RECT 5.86 1.12 6.18 1.4 ;
  LAYER M3 ;
        RECT 5.88 1.1 6.16 1.42 ;
  LAYER M2 ;
        RECT 6.72 1.12 7.04 1.4 ;
  LAYER M3 ;
        RECT 6.74 1.1 7.02 1.42 ;
  LAYER M2 ;
        RECT 5.86 0.7 6.18 0.98 ;
  LAYER M3 ;
        RECT 5.88 0.68 6.16 1 ;
  LAYER M2 ;
        RECT 5.86 1.12 6.18 1.4 ;
  LAYER M3 ;
        RECT 5.88 1.1 6.16 1.42 ;
  LAYER M2 ;
        RECT 6.72 1.12 7.04 1.4 ;
  LAYER M3 ;
        RECT 6.74 1.1 7.02 1.42 ;
  LAYER M2 ;
        RECT 5.86 0.7 6.18 0.98 ;
  LAYER M3 ;
        RECT 5.88 0.68 6.16 1 ;
  LAYER M2 ;
        RECT 5.86 1.12 6.18 1.4 ;
  LAYER M3 ;
        RECT 5.88 1.1 6.16 1.42 ;
  LAYER M2 ;
        RECT 6.72 1.12 7.04 1.4 ;
  LAYER M3 ;
        RECT 6.74 1.1 7.02 1.42 ;
  LAYER M2 ;
        RECT 0.26 2.8 1.46 3.08 ;
  LAYER M2 ;
        RECT 0.26 12.04 1.46 12.32 ;
  LAYER M2 ;
        RECT 0.27 2.8 0.59 3.08 ;
  LAYER M3 ;
        RECT 0.29 2.94 0.57 12.18 ;
  LAYER M2 ;
        RECT 0.27 12.04 0.59 12.32 ;
  LAYER M2 ;
        RECT 2.84 10.36 4.04 10.64 ;
  LAYER M3 ;
        RECT 0.29 10.315 0.57 10.685 ;
  LAYER M2 ;
        RECT 0.43 10.36 3.01 10.64 ;
  LAYER M2 ;
        RECT 0.27 10.36 0.59 10.64 ;
  LAYER M3 ;
        RECT 0.29 10.34 0.57 10.66 ;
  LAYER M2 ;
        RECT 0.27 10.36 0.59 10.64 ;
  LAYER M3 ;
        RECT 0.29 10.34 0.57 10.66 ;
  LAYER M2 ;
        RECT 7.14 2.8 8.34 3.08 ;
  LAYER M2 ;
        RECT 9.72 2.8 10.92 3.08 ;
  LAYER M2 ;
        RECT 9.72 12.04 10.92 12.32 ;
  LAYER M2 ;
        RECT 9.73 2.8 10.05 3.08 ;
  LAYER M3 ;
        RECT 9.75 2.94 10.03 12.18 ;
  LAYER M2 ;
        RECT 9.73 12.04 10.05 12.32 ;
  LAYER M2 ;
        RECT 8.17 2.8 9.89 3.08 ;
  LAYER M2 ;
        RECT 2.84 14.56 4.04 14.84 ;
  LAYER M3 ;
        RECT 2.44 15.38 2.72 19.9 ;
  LAYER M2 ;
        RECT 2.58 14.56 3.01 14.84 ;
  LAYER M3 ;
        RECT 2.44 14.7 2.72 15.54 ;
  LAYER M2 ;
        RECT 2.42 14.56 2.74 14.84 ;
  LAYER M3 ;
        RECT 2.44 14.54 2.72 14.86 ;
  LAYER M2 ;
        RECT 2.42 14.56 2.74 14.84 ;
  LAYER M3 ;
        RECT 2.44 14.54 2.72 14.86 ;
  LAYER M2 ;
        RECT 7.14 14.56 8.34 14.84 ;
  LAYER M3 ;
        RECT 8.46 15.38 8.74 19.9 ;
  LAYER M2 ;
        RECT 8.17 14.56 8.6 14.84 ;
  LAYER M3 ;
        RECT 8.46 14.7 8.74 15.54 ;
  LAYER M2 ;
        RECT 8.44 14.56 8.76 14.84 ;
  LAYER M3 ;
        RECT 8.46 14.54 8.74 14.86 ;
  LAYER M2 ;
        RECT 8.44 14.56 8.76 14.84 ;
  LAYER M3 ;
        RECT 8.46 14.54 8.74 14.86 ;
  LAYER M1 ;
        RECT 5.895 15.455 6.145 18.985 ;
  LAYER M1 ;
        RECT 5.895 19.235 6.145 20.245 ;
  LAYER M1 ;
        RECT 5.895 21.335 6.145 22.345 ;
  LAYER M1 ;
        RECT 6.325 15.455 6.575 18.985 ;
  LAYER M1 ;
        RECT 5.465 15.455 5.715 18.985 ;
  LAYER M1 ;
        RECT 5.035 15.455 5.285 18.985 ;
  LAYER M1 ;
        RECT 5.035 19.235 5.285 20.245 ;
  LAYER M1 ;
        RECT 5.035 21.335 5.285 22.345 ;
  LAYER M1 ;
        RECT 4.605 15.455 4.855 18.985 ;
  LAYER M2 ;
        RECT 5.85 15.4 7.05 15.68 ;
  LAYER M2 ;
        RECT 4.99 19.6 6.19 19.88 ;
  LAYER M2 ;
        RECT 4.99 21.7 6.19 21.98 ;
  LAYER M2 ;
        RECT 4.56 16.24 6.62 16.52 ;
  LAYER M3 ;
        RECT 5.88 15.38 6.16 19.9 ;
  LAYER M2 ;
        RECT 4.99 15.82 6.19 16.1 ;
  LAYER M3 ;
        RECT 5.02 16.22 5.3 22 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 3.865 ;
  LAYER M1 ;
        RECT 3.745 4.115 3.995 5.125 ;
  LAYER M1 ;
        RECT 3.745 6.215 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.315 0.335 3.565 3.865 ;
  LAYER M1 ;
        RECT 4.175 0.335 4.425 3.865 ;
  LAYER M1 ;
        RECT 4.605 0.335 4.855 3.865 ;
  LAYER M1 ;
        RECT 4.605 4.115 4.855 5.125 ;
  LAYER M1 ;
        RECT 4.605 6.215 4.855 7.225 ;
  LAYER M1 ;
        RECT 5.035 0.335 5.285 3.865 ;
  LAYER M2 ;
        RECT 2.84 0.28 4.04 0.56 ;
  LAYER M2 ;
        RECT 3.7 4.48 4.9 4.76 ;
  LAYER M2 ;
        RECT 3.7 6.58 4.9 6.86 ;
  LAYER M2 ;
        RECT 3.27 1.12 5.33 1.4 ;
  LAYER M3 ;
        RECT 3.73 0.26 4.01 4.78 ;
  LAYER M2 ;
        RECT 3.7 0.7 4.9 0.98 ;
  LAYER M3 ;
        RECT 4.59 1.1 4.87 6.88 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 14.785 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M2 ;
        RECT 0.69 8.26 1.89 8.54 ;
  LAYER M2 ;
        RECT 0.69 14.14 1.89 14.42 ;
  LAYER M2 ;
        RECT 0.26 7.84 1.46 8.12 ;
  LAYER M2 ;
        RECT 0.26 12.04 1.46 12.32 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 14.44 ;
  LAYER M1 ;
        RECT 1.165 3.695 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.165 2.435 1.415 3.445 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 1.345 ;
  LAYER M1 ;
        RECT 0.735 3.695 0.985 7.225 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M2 ;
        RECT 0.69 6.58 1.89 6.86 ;
  LAYER M2 ;
        RECT 0.69 0.7 1.89 0.98 ;
  LAYER M2 ;
        RECT 0.26 7 1.46 7.28 ;
  LAYER M2 ;
        RECT 0.26 2.8 1.46 3.08 ;
  LAYER M3 ;
        RECT 1.58 0.68 1.86 6.88 ;
  LAYER M1 ;
        RECT 9.765 7.895 10.015 11.425 ;
  LAYER M1 ;
        RECT 9.765 11.675 10.015 12.685 ;
  LAYER M1 ;
        RECT 9.765 13.775 10.015 14.785 ;
  LAYER M1 ;
        RECT 10.195 7.895 10.445 11.425 ;
  LAYER M1 ;
        RECT 9.335 7.895 9.585 11.425 ;
  LAYER M2 ;
        RECT 9.29 8.26 10.49 8.54 ;
  LAYER M2 ;
        RECT 9.29 14.14 10.49 14.42 ;
  LAYER M2 ;
        RECT 9.72 7.84 10.92 8.12 ;
  LAYER M2 ;
        RECT 9.72 12.04 10.92 12.32 ;
  LAYER M3 ;
        RECT 9.32 8.24 9.6 14.44 ;
  LAYER M1 ;
        RECT 9.765 3.695 10.015 7.225 ;
  LAYER M1 ;
        RECT 9.765 2.435 10.015 3.445 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 1.345 ;
  LAYER M1 ;
        RECT 10.195 3.695 10.445 7.225 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M2 ;
        RECT 9.29 6.58 10.49 6.86 ;
  LAYER M2 ;
        RECT 9.29 0.7 10.49 0.98 ;
  LAYER M2 ;
        RECT 9.72 7 10.92 7.28 ;
  LAYER M2 ;
        RECT 9.72 2.8 10.92 3.08 ;
  LAYER M3 ;
        RECT 9.32 0.68 9.6 6.88 ;
  LAYER M1 ;
        RECT 3.745 11.255 3.995 14.785 ;
  LAYER M1 ;
        RECT 3.745 9.995 3.995 11.005 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 8.905 ;
  LAYER M1 ;
        RECT 3.315 11.255 3.565 14.785 ;
  LAYER M1 ;
        RECT 4.175 11.255 4.425 14.785 ;
  LAYER M1 ;
        RECT 4.605 11.255 4.855 14.785 ;
  LAYER M1 ;
        RECT 4.605 9.995 4.855 11.005 ;
  LAYER M1 ;
        RECT 4.605 7.895 4.855 8.905 ;
  LAYER M1 ;
        RECT 5.035 11.255 5.285 14.785 ;
  LAYER M2 ;
        RECT 3.7 8.26 5.33 8.54 ;
  LAYER M2 ;
        RECT 3.27 13.72 5.33 14 ;
  LAYER M2 ;
        RECT 2.84 14.56 4.04 14.84 ;
  LAYER M2 ;
        RECT 3.7 14.14 4.9 14.42 ;
  LAYER M2 ;
        RECT 2.84 10.36 4.04 10.64 ;
  LAYER M2 ;
        RECT 3.7 9.94 4.9 10.22 ;
  LAYER M3 ;
        RECT 5.02 8.24 5.3 14.02 ;
  LAYER M1 ;
        RECT 8.475 15.455 8.725 18.985 ;
  LAYER M1 ;
        RECT 8.475 19.235 8.725 20.245 ;
  LAYER M1 ;
        RECT 8.475 21.335 8.725 22.345 ;
  LAYER M1 ;
        RECT 8.905 15.455 9.155 18.985 ;
  LAYER M1 ;
        RECT 8.045 15.455 8.295 18.985 ;
  LAYER M2 ;
        RECT 8.43 15.4 9.63 15.68 ;
  LAYER M2 ;
        RECT 8.43 19.6 9.63 19.88 ;
  LAYER M2 ;
        RECT 8 15.82 9.2 16.1 ;
  LAYER M2 ;
        RECT 8 21.7 9.2 21.98 ;
  LAYER M3 ;
        RECT 8.46 15.38 8.74 19.9 ;
  LAYER M3 ;
        RECT 8.03 15.8 8.31 22 ;
  LAYER M1 ;
        RECT 2.455 15.455 2.705 18.985 ;
  LAYER M1 ;
        RECT 2.455 19.235 2.705 20.245 ;
  LAYER M1 ;
        RECT 2.455 21.335 2.705 22.345 ;
  LAYER M1 ;
        RECT 2.025 15.455 2.275 18.985 ;
  LAYER M1 ;
        RECT 2.885 15.455 3.135 18.985 ;
  LAYER M2 ;
        RECT 1.55 15.4 2.75 15.68 ;
  LAYER M2 ;
        RECT 1.55 19.6 2.75 19.88 ;
  LAYER M2 ;
        RECT 1.98 15.82 3.18 16.1 ;
  LAYER M2 ;
        RECT 1.98 21.7 3.18 21.98 ;
  LAYER M3 ;
        RECT 2.44 15.38 2.72 19.9 ;
  LAYER M3 ;
        RECT 2.87 15.8 3.15 22 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.185 2.435 7.435 3.445 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 1.345 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M2 ;
        RECT 6.71 6.58 7.91 6.86 ;
  LAYER M2 ;
        RECT 6.71 0.7 7.91 0.98 ;
  LAYER M2 ;
        RECT 7.14 7 8.34 7.28 ;
  LAYER M2 ;
        RECT 7.14 2.8 8.34 3.08 ;
  LAYER M3 ;
        RECT 6.74 0.68 7.02 6.88 ;
  LAYER M1 ;
        RECT 7.185 11.255 7.435 14.785 ;
  LAYER M1 ;
        RECT 7.185 9.995 7.435 11.005 ;
  LAYER M1 ;
        RECT 7.185 7.895 7.435 8.905 ;
  LAYER M1 ;
        RECT 7.615 11.255 7.865 14.785 ;
  LAYER M1 ;
        RECT 6.755 11.255 7.005 14.785 ;
  LAYER M2 ;
        RECT 6.71 14.14 7.91 14.42 ;
  LAYER M2 ;
        RECT 6.71 8.26 7.91 8.54 ;
  LAYER M2 ;
        RECT 7.14 14.56 8.34 14.84 ;
  LAYER M2 ;
        RECT 7.14 10.36 8.34 10.64 ;
  LAYER M3 ;
        RECT 6.74 8.24 7.02 14.44 ;
  END 
END CP
