MACRO TELESCOPIC_OTA
  ORIGIN 0 0 ;
  FOREIGN TELESCOPIC_OTA 0 0 ;
  SIZE 1.492 BY 11.844 ;
  PIN ID
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 0.3 1.392 0.34 2.304 ;
    END
  END ID
  PIN VBIASP2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.444 10.316 0.996 10.348 ;
    END
  END VBIASP2
  PIN VOUTN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.844 6.956 1.076 6.988 ;
      LAYER M2 ;
        RECT 0.844 7.124 1.076 7.156 ;
      LAYER M2 ;
        RECT 0.844 6.956 0.916 6.988 ;
      LAYER M1 ;
        RECT 0.864 6.966 0.896 7.146 ;
      LAYER M2 ;
        RECT 0.844 7.124 0.916 7.156 ;
    END
  END VOUTN
  PIN VOUTP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.364 6.872 0.596 6.904 ;
      LAYER M2 ;
        RECT 0.364 7.208 0.596 7.24 ;
      LAYER M2 ;
        RECT 0.524 6.872 0.596 6.904 ;
      LAYER M1 ;
        RECT 0.544 6.888 0.576 7.224 ;
      LAYER M2 ;
        RECT 0.524 7.208 0.596 7.24 ;
    END
  END VOUTP
  PIN VBIASN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.364 6.116 1.076 6.148 ;
    END
  END VBIASN
  PIN VBIASP1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.364 7.964 1.076 7.996 ;
    END
  END VBIASP1
  PIN VINP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.444 3.764 1.156 3.796 ;
    END
  END VINP
  PIN VINN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.284 3.68 0.996 3.712 ;
    END
  END VINN
  OBS 
  LAYER M2 ;
        RECT 0.444 2.168 0.676 2.2 ;
  LAYER M2 ;
        RECT 0.204 4.436 1.236 4.468 ;
  LAYER M2 ;
        RECT 0.524 2.168 0.596 2.2 ;
  LAYER M3 ;
        RECT 0.54 2.184 0.58 4.452 ;
  LAYER M2 ;
        RECT 0.524 4.436 0.596 4.468 ;
  LAYER M2 ;
        RECT 0.524 2.168 0.596 2.2 ;
  LAYER M3 ;
        RECT 0.54 2.148 0.58 2.22 ;
  LAYER M2 ;
        RECT 0.524 4.436 0.596 4.468 ;
  LAYER M3 ;
        RECT 0.54 4.416 0.58 4.488 ;
  LAYER M2 ;
        RECT 0.524 2.168 0.596 2.2 ;
  LAYER M3 ;
        RECT 0.54 2.148 0.58 2.22 ;
  LAYER M2 ;
        RECT 0.524 4.436 0.596 4.468 ;
  LAYER M3 ;
        RECT 0.54 4.416 0.58 4.488 ;
  LAYER M2 ;
        RECT 0.284 7.376 0.516 7.408 ;
  LAYER M2 ;
        RECT 0.444 9.476 0.996 9.508 ;
  LAYER M2 ;
        RECT 0.444 7.376 0.516 7.408 ;
  LAYER M3 ;
        RECT 0.46 7.392 0.5 9.492 ;
  LAYER M2 ;
        RECT 0.444 9.476 0.516 9.508 ;
  LAYER M2 ;
        RECT 0.444 7.376 0.516 7.408 ;
  LAYER M3 ;
        RECT 0.46 7.356 0.5 7.428 ;
  LAYER M2 ;
        RECT 0.444 9.476 0.516 9.508 ;
  LAYER M3 ;
        RECT 0.46 9.456 0.5 9.528 ;
  LAYER M2 ;
        RECT 0.444 7.376 0.516 7.408 ;
  LAYER M3 ;
        RECT 0.46 7.356 0.5 7.428 ;
  LAYER M2 ;
        RECT 0.444 9.476 0.516 9.508 ;
  LAYER M3 ;
        RECT 0.46 9.456 0.5 9.528 ;
  LAYER M2 ;
        RECT 0.924 7.292 1.156 7.324 ;
  LAYER M2 ;
        RECT 0.604 9.56 0.836 9.592 ;
  LAYER M2 ;
        RECT 0.8 7.292 0.96 7.324 ;
  LAYER M3 ;
        RECT 0.78 7.308 0.82 9.576 ;
  LAYER M2 ;
        RECT 0.764 9.56 0.836 9.592 ;
  LAYER M2 ;
        RECT 0.764 7.292 0.836 7.324 ;
  LAYER M3 ;
        RECT 0.78 7.272 0.82 7.344 ;
  LAYER M2 ;
        RECT 0.764 9.56 0.836 9.592 ;
  LAYER M3 ;
        RECT 0.78 9.54 0.82 9.612 ;
  LAYER M2 ;
        RECT 0.764 7.292 0.836 7.324 ;
  LAYER M3 ;
        RECT 0.78 7.272 0.82 7.344 ;
  LAYER M2 ;
        RECT 0.764 9.56 0.836 9.592 ;
  LAYER M3 ;
        RECT 0.78 9.54 0.82 9.612 ;
  LAYER M2 ;
        RECT 0.444 4.604 1.156 4.636 ;
  LAYER M2 ;
        RECT 0.924 6.788 1.156 6.82 ;
  LAYER M2 ;
        RECT 0.924 4.604 0.996 4.636 ;
  LAYER M3 ;
        RECT 0.94 4.62 0.98 6.804 ;
  LAYER M2 ;
        RECT 0.924 6.788 0.996 6.82 ;
  LAYER M2 ;
        RECT 0.924 4.604 0.996 4.636 ;
  LAYER M3 ;
        RECT 0.94 4.584 0.98 4.656 ;
  LAYER M2 ;
        RECT 0.924 6.788 0.996 6.82 ;
  LAYER M3 ;
        RECT 0.94 6.768 0.98 6.84 ;
  LAYER M2 ;
        RECT 0.924 4.604 0.996 4.636 ;
  LAYER M3 ;
        RECT 0.94 4.584 0.98 4.656 ;
  LAYER M2 ;
        RECT 0.924 6.788 0.996 6.82 ;
  LAYER M3 ;
        RECT 0.94 6.768 0.98 6.84 ;
  LAYER M2 ;
        RECT 0.284 4.52 0.996 4.552 ;
  LAYER M2 ;
        RECT 0.284 6.704 0.516 6.736 ;
  LAYER M2 ;
        RECT 0.284 4.52 0.356 4.552 ;
  LAYER M3 ;
        RECT 0.3 4.536 0.34 6.72 ;
  LAYER M2 ;
        RECT 0.284 6.704 0.356 6.736 ;
  LAYER M2 ;
        RECT 0.284 4.52 0.356 4.552 ;
  LAYER M3 ;
        RECT 0.3 4.5 0.34 4.572 ;
  LAYER M2 ;
        RECT 0.284 6.704 0.356 6.736 ;
  LAYER M3 ;
        RECT 0.3 6.684 0.34 6.756 ;
  LAYER M2 ;
        RECT 0.284 4.52 0.356 4.552 ;
  LAYER M3 ;
        RECT 0.3 4.5 0.34 4.572 ;
  LAYER M2 ;
        RECT 0.284 6.704 0.356 6.736 ;
  LAYER M3 ;
        RECT 0.3 6.684 0.34 6.756 ;
  LAYER M1 ;
        RECT 0.304 1.56 0.336 2.304 ;
  LAYER M1 ;
        RECT 0.304 1.224 0.336 1.464 ;
  LAYER M1 ;
        RECT 0.304 0.468 0.336 0.708 ;
  LAYER M1 ;
        RECT 0.224 1.56 0.256 2.304 ;
  LAYER M1 ;
        RECT 0.384 1.56 0.416 2.304 ;
  LAYER M1 ;
        RECT 0.464 1.56 0.496 2.304 ;
  LAYER M1 ;
        RECT 0.464 1.224 0.496 1.464 ;
  LAYER M1 ;
        RECT 0.464 0.468 0.496 0.708 ;
  LAYER M1 ;
        RECT 0.544 1.56 0.576 2.304 ;
  LAYER M1 ;
        RECT 0.624 1.56 0.656 2.304 ;
  LAYER M1 ;
        RECT 0.624 1.224 0.656 1.464 ;
  LAYER M1 ;
        RECT 0.624 0.468 0.656 0.708 ;
  LAYER M1 ;
        RECT 0.704 1.56 0.736 2.304 ;
  LAYER M1 ;
        RECT 0.784 1.56 0.816 2.304 ;
  LAYER M1 ;
        RECT 0.784 1.224 0.816 1.464 ;
  LAYER M1 ;
        RECT 0.784 0.468 0.816 0.708 ;
  LAYER M1 ;
        RECT 0.864 1.56 0.896 2.304 ;
  LAYER M2 ;
        RECT 0.284 2.252 0.836 2.284 ;
  LAYER M2 ;
        RECT 0.284 1.412 0.836 1.444 ;
  LAYER M2 ;
        RECT 0.204 2.084 0.916 2.116 ;
  LAYER M2 ;
        RECT 0.284 0.572 0.836 0.604 ;
  LAYER M3 ;
        RECT 0.3 1.392 0.34 2.304 ;
  LAYER M2 ;
        RECT 0.444 2.168 0.676 2.2 ;
  LAYER M3 ;
        RECT 0.46 0.552 0.5 2.136 ;
  LAYER M1 ;
        RECT 0.464 9.456 0.496 10.2 ;
  LAYER M1 ;
        RECT 0.464 10.296 0.496 10.536 ;
  LAYER M1 ;
        RECT 0.464 11.052 0.496 11.292 ;
  LAYER M1 ;
        RECT 0.384 9.456 0.416 10.2 ;
  LAYER M1 ;
        RECT 0.544 9.456 0.576 10.2 ;
  LAYER M1 ;
        RECT 0.624 9.456 0.656 10.2 ;
  LAYER M1 ;
        RECT 0.624 10.296 0.656 10.536 ;
  LAYER M1 ;
        RECT 0.624 11.052 0.656 11.292 ;
  LAYER M1 ;
        RECT 0.704 9.456 0.736 10.2 ;
  LAYER M1 ;
        RECT 0.784 9.456 0.816 10.2 ;
  LAYER M1 ;
        RECT 0.784 10.296 0.816 10.536 ;
  LAYER M1 ;
        RECT 0.784 11.052 0.816 11.292 ;
  LAYER M1 ;
        RECT 0.864 9.456 0.896 10.2 ;
  LAYER M1 ;
        RECT 0.944 9.456 0.976 10.2 ;
  LAYER M1 ;
        RECT 0.944 10.296 0.976 10.536 ;
  LAYER M1 ;
        RECT 0.944 11.052 0.976 11.292 ;
  LAYER M1 ;
        RECT 1.024 9.456 1.056 10.2 ;
  LAYER M2 ;
        RECT 0.364 9.644 1.076 9.676 ;
  LAYER M2 ;
        RECT 0.444 11.156 0.996 11.188 ;
  LAYER M2 ;
        RECT 0.444 9.476 0.996 9.508 ;
  LAYER M2 ;
        RECT 0.604 9.56 0.836 9.592 ;
  LAYER M2 ;
        RECT 0.444 10.316 0.996 10.348 ;
  LAYER M3 ;
        RECT 0.7 9.624 0.74 11.208 ;
  LAYER M1 ;
        RECT 1.024 6.264 1.056 7.008 ;
  LAYER M1 ;
        RECT 1.024 5.928 1.056 6.168 ;
  LAYER M1 ;
        RECT 1.024 5.172 1.056 5.412 ;
  LAYER M1 ;
        RECT 1.104 6.264 1.136 7.008 ;
  LAYER M1 ;
        RECT 0.944 6.264 0.976 7.008 ;
  LAYER M1 ;
        RECT 0.384 6.264 0.416 7.008 ;
  LAYER M1 ;
        RECT 0.384 5.928 0.416 6.168 ;
  LAYER M1 ;
        RECT 0.384 5.172 0.416 5.412 ;
  LAYER M1 ;
        RECT 0.464 6.264 0.496 7.008 ;
  LAYER M1 ;
        RECT 0.304 6.264 0.336 7.008 ;
  LAYER M2 ;
        RECT 0.364 5.276 1.076 5.308 ;
  LAYER M2 ;
        RECT 0.844 6.956 1.076 6.988 ;
  LAYER M2 ;
        RECT 0.364 6.872 0.596 6.904 ;
  LAYER M2 ;
        RECT 0.364 6.116 1.076 6.148 ;
  LAYER M2 ;
        RECT 0.924 6.788 1.156 6.82 ;
  LAYER M2 ;
        RECT 0.284 6.704 0.516 6.736 ;
  LAYER M1 ;
        RECT 1.024 7.104 1.056 7.848 ;
  LAYER M1 ;
        RECT 1.024 7.944 1.056 8.184 ;
  LAYER M1 ;
        RECT 1.024 8.7 1.056 8.94 ;
  LAYER M1 ;
        RECT 1.104 7.104 1.136 7.848 ;
  LAYER M1 ;
        RECT 0.944 7.104 0.976 7.848 ;
  LAYER M1 ;
        RECT 0.384 7.104 0.416 7.848 ;
  LAYER M1 ;
        RECT 0.384 7.944 0.416 8.184 ;
  LAYER M1 ;
        RECT 0.384 8.7 0.416 8.94 ;
  LAYER M1 ;
        RECT 0.464 7.104 0.496 7.848 ;
  LAYER M1 ;
        RECT 0.304 7.104 0.336 7.848 ;
  LAYER M2 ;
        RECT 0.364 8.804 1.076 8.836 ;
  LAYER M2 ;
        RECT 0.844 7.124 1.076 7.156 ;
  LAYER M2 ;
        RECT 0.364 7.208 0.596 7.24 ;
  LAYER M2 ;
        RECT 0.364 7.964 1.076 7.996 ;
  LAYER M2 ;
        RECT 0.924 7.292 1.156 7.324 ;
  LAYER M2 ;
        RECT 0.284 7.376 0.516 7.408 ;
  LAYER M1 ;
        RECT 1.104 3.912 1.136 4.656 ;
  LAYER M1 ;
        RECT 1.104 3.576 1.136 3.816 ;
  LAYER M1 ;
        RECT 1.104 2.82 1.136 3.06 ;
  LAYER M1 ;
        RECT 1.184 3.912 1.216 4.656 ;
  LAYER M1 ;
        RECT 1.024 3.912 1.056 4.656 ;
  LAYER M1 ;
        RECT 0.944 3.912 0.976 4.656 ;
  LAYER M1 ;
        RECT 0.944 3.576 0.976 3.816 ;
  LAYER M1 ;
        RECT 0.944 2.82 0.976 3.06 ;
  LAYER M1 ;
        RECT 0.864 3.912 0.896 4.656 ;
  LAYER M1 ;
        RECT 0.784 3.912 0.816 4.656 ;
  LAYER M1 ;
        RECT 0.784 3.576 0.816 3.816 ;
  LAYER M1 ;
        RECT 0.784 2.82 0.816 3.06 ;
  LAYER M1 ;
        RECT 0.704 3.912 0.736 4.656 ;
  LAYER M1 ;
        RECT 0.624 3.912 0.656 4.656 ;
  LAYER M1 ;
        RECT 0.624 3.576 0.656 3.816 ;
  LAYER M1 ;
        RECT 0.624 2.82 0.656 3.06 ;
  LAYER M1 ;
        RECT 0.544 3.912 0.576 4.656 ;
  LAYER M1 ;
        RECT 0.464 3.912 0.496 4.656 ;
  LAYER M1 ;
        RECT 0.464 3.576 0.496 3.816 ;
  LAYER M1 ;
        RECT 0.464 2.82 0.496 3.06 ;
  LAYER M1 ;
        RECT 0.384 3.912 0.416 4.656 ;
  LAYER M1 ;
        RECT 0.304 3.912 0.336 4.656 ;
  LAYER M1 ;
        RECT 0.304 3.576 0.336 3.816 ;
  LAYER M1 ;
        RECT 0.304 2.82 0.336 3.06 ;
  LAYER M1 ;
        RECT 0.224 3.912 0.256 4.656 ;
  LAYER M2 ;
        RECT 0.284 2.924 1.156 2.956 ;
  LAYER M2 ;
        RECT 0.444 4.604 1.156 4.636 ;
  LAYER M2 ;
        RECT 0.284 4.52 0.996 4.552 ;
  LAYER M2 ;
        RECT 0.444 3.764 1.156 3.796 ;
  LAYER M2 ;
        RECT 0.284 3.68 0.996 3.712 ;
  LAYER M2 ;
        RECT 0.204 4.436 1.236 4.468 ;
  END 
END TELESCOPIC_OTA
